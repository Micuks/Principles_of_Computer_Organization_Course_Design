module cpu (
    input clr,
    input t3,
    input swa,
    input swb,
    input swc,
    input ir4,
    input ir5,
    input ir6,
    input ir7,
    input w1,
    input w2,
    input w3,
    input c,
    input z,
    output drw,
    output pcinc,
    output lpc,
    output lar,
    output pcadd,
    output arinc,
    output selctl,
    output memw,
    output stop,
    output lir,
    output ldz,
    output ldc,
    output cin,
    output s0,
    output s1,
    output s2,
    output s3,
    output m,
    output abus,
    output sbus,
    output mbus,
    output short,
    output long,
    output sel0,
    output sel1,
    output sel2,
    output sel3);
    
endmodule